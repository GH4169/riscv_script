wildcard vadd.vv = {32'b000000_?_?????_?????_000_?????_1010111};
wildcard vadd.vx = {32'b000000_?_?????_?????_100_?????_1010111};
wildcard vadd.vi = {32'b000000_?_?????_?????_011_?????_1010111};
wildcard vsub.vv = {32'b000010_?_?????_?????_000_?????_1010111};
wildcard vsub.vx = {32'b000010_?_?????_?????_100_?????_1010111};
wildcard vrsub.vx = {32'b000011_?_?????_?????_100_?????_1010111};
wildcard vrsub.vi = {32'b000011_?_?????_?????_011_?????_1010111};
wildcard vwaddu.vv = {32'b110000_?_?????_?????_010_?????_1010111};
wildcard vwaddu.vx = {32'b110000_?_?????_?????_110_?????_1010111};
wildcard vwsubu.vv = {32'b110010_?_?????_?????_010_?????_1010111};
wildcard vwsubu.vx = {32'b110010_?_?????_?????_110_?????_1010111};
wildcard vwadd.vv = {32'b110001_?_?????_?????_010_?????_1010111};
wildcard vwadd.vx = {32'b110001_?_?????_?????_110_?????_1010111};
wildcard vwsub.vv = {32'b110011_?_?????_?????_010_?????_1010111};
wildcard vwsub.vx = {32'b110011_?_?????_?????_110_?????_1010111};
wildcard vwaddu.wv = {32'b110100_?_?????_?????_010_?????_1010111};
wildcard vwaddu.wx = {32'b110100_?_?????_?????_110_?????_1010111};
wildcard vwsubu.wv = {32'b110110_?_?????_?????_010_?????_1010111};
wildcard vwsubu.wx = {32'b110110_?_?????_?????_110_?????_1010111};
wildcard vwadd.wv = {32'b110101_?_?????_?????_010_?????_1010111};
wildcard vwadd.wx = {32'b110101_?_?????_?????_110_?????_1010111};
wildcard vwsub.wv = {32'b110111_?_?????_?????_010_?????_1010111};
wildcard vwsub.wx = {32'b110111_?_?????_?????_110_?????_1010111};
wildcard vzext.vf2 = {32'b010010_?_?????_00110_010_?????_1010111};
wildcard vsext.vf2 = {32'b010010_?_?????_00111_010_?????_1010111};
wildcard vzext.vf4 = {32'b010010_?_?????_00100_010_?????_1010111};
wildcard vsext.vf4 = {32'b010010_?_?????_00101_010_?????_1010111};
wildcard vzext.vf8 = {32'b010010_?_?????_00010_010_?????_1010111};
wildcard vsext.vf8 = {32'b010010_?_?????_00011_010_?????_1010111};
wildcard vadc.vvm = {32'b010000_0_?????_?????_000_?????_1010111};
wildcard vadc.vxm = {32'b010000_0_?????_?????_100_?????_1010111};
wildcard vadc.vim = {32'b010000_0_?????_?????_011_?????_1010111};
wildcard vmadc.vvm = {32'b010001_0_?????_?????_000_?????_1010111};
wildcard vmadc.vxm = {32'b010001_0_?????_?????_100_?????_1010111};
wildcard vmadc.vim = {32'b010001_0_?????_?????_011_?????_1010111};
wildcard vmadc.vv = {32'b010001_1_?????_?????_000_?????_1010111};
wildcard vmadc.vx = {32'b010001_1_?????_?????_100_?????_1010111};
wildcard vmadc.vi = {32'b010001_1_?????_?????_011_?????_1010111};
wildcard vsbc.vvm = {32'b010010_0_?????_?????_000_?????_1010111};
wildcard vsbc.vxm = {32'b010010_0_?????_?????_100_?????_1010111};
wildcard vmsbc.vvm = {32'b010011_0_?????_?????_000_?????_1010111};
wildcard vmsbc.vxm = {32'b010011_0_?????_?????_100_?????_1010111};
wildcard vmsbc.vv = {32'b010011_1_?????_?????_000_?????_1010111};
wildcard vmsbc.vx = {32'b010011_1_?????_?????_100_?????_1010111};
wildcard vand.vv = {32'b001001_?_?????_?????_000_?????_1010111};
wildcard vand.vx = {32'b001001_?_?????_?????_100_?????_1010111};
wildcard vand.vi = {32'b001001_?_?????_?????_011_?????_1010111};
wildcard vor.vv = {32'b001010_?_?????_?????_000_?????_1010111};
wildcard vor.vx = {32'b001010_?_?????_?????_100_?????_1010111};
wildcard vor.vi = {32'b001010_?_?????_?????_011_?????_1010111};
wildcard vxor.vv = {32'b001011_?_?????_?????_000_?????_1010111};
wildcard vxor.vx = {32'b001011_?_?????_?????_100_?????_1010111};
wildcard vxor.vi = {32'b001011_?_?????_?????_011_?????_1010111};
wildcard vsll.vv = {32'b100101_?_?????_?????_000_?????_1010111};
wildcard vsll.vx = {32'b100101_?_?????_?????_100_?????_1010111};
wildcard vsll.vi = {32'b100101_?_?????_?????_011_?????_1010111};
wildcard vsrl.vv = {32'b101000_?_?????_?????_000_?????_1010111};
wildcard vsrl.vx = {32'b101000_?_?????_?????_100_?????_1010111};
wildcard vsrl.vi = {32'b101000_?_?????_?????_011_?????_1010111};
wildcard vsra.vv = {32'b101001_?_?????_?????_000_?????_1010111};
wildcard vsra.vx = {32'b101001_?_?????_?????_100_?????_1010111};
wildcard vsra.vi = {32'b101001_?_?????_?????_011_?????_1010111};
wildcard vnsrl.wv = {32'b101100_?_?????_?????_000_?????_1010111};
wildcard vnsrl.wx = {32'b101100_?_?????_?????_100_?????_1010111};
wildcard vnsrl.wi = {32'b101100_?_?????_?????_011_?????_1010111};
wildcard vnsra.wv = {32'b101101_?_?????_?????_000_?????_1010111};
wildcard vnsra.wx = {32'b101101_?_?????_?????_100_?????_1010111};
wildcard vnsra.wi = {32'b101101_?_?????_?????_011_?????_1010111};
wildcard vmseq.vv = {32'b011000_?_?????_?????_000_?????_1010111};
wildcard vmseq.vx = {32'b011000_?_?????_?????_100_?????_1010111};
wildcard vmseq.vi = {32'b011000_?_?????_?????_011_?????_1010111};
wildcard vmsne.vv = {32'b011001_?_?????_?????_000_?????_1010111};
wildcard vmsne.vx = {32'b011001_?_?????_?????_100_?????_1010111};
wildcard vmsne.vi = {32'b011001_?_?????_?????_011_?????_1010111};
wildcard vmsltu.vv = {32'b011010_?_?????_?????_000_?????_1010111};
wildcard vmsltu.vx = {32'b011010_?_?????_?????_100_?????_1010111};
wildcard vmslt.vv = {32'b011011_?_?????_?????_000_?????_1010111};
wildcard vmslt.vx = {32'b011011_?_?????_?????_100_?????_1010111};
wildcard vmsleu.vv = {32'b11100_?_?????_?????_000_?????_1010111};
wildcard vmsleu.vx = {32'b11100_?_?????_?????_100_?????_1010111};
wildcard vmsleu.vi = {32'b11100_?_?????_?????_011_?????_1010111};
wildcard vmsle.vv = {32'b011101_?_?????_?????_000_?????_1010111};
wildcard vmsle.vx = {32'b011101_?_?????_?????_100_?????_1010111};
wildcard vmsle.vi = {32'b011101_?_?????_?????_011_?????_1010111};
wildcard vmsgtu.vx = {32'b011110_?_?????_?????_100_?????_1010111};
wildcard vmsgtu.vi = {32'b011110_?_?????_?????_011_?????_1010111};
wildcard vmsgt.vx = {32'b011111_?_?????_?????_100_?????_1010111};
wildcard vmsgt.vi = {32'b011111_?_?????_?????_011_?????_1010111};
wildcard vminu.vv = {32'b000100_?_?????_?????_000_?????_1010111};
wildcard vminu.vx = {32'b000100_?_?????_?????_100_?????_1010111};
wildcard vmin.vv = {32'b000101_?_?????_?????_000_?????_1010111};
wildcard vmin.vx = {32'b000101_?_?????_?????_100_?????_1010111};
wildcard vmaxu.vv = {32'b000110_?_?????_?????_000_?????_1010111};
wildcard vmaxu.vx = {32'b000110_?_?????_?????_100_?????_1010111};
wildcard vmax.vv = {32'b000111_?_?????_?????_000_?????_1010111};
wildcard vmax.vx = {32'b000111_?_?????_?????_100_?????_1010111};
wildcard vmul.vv = {32'b100101_?_?????_?????_010_?????_1010111};
wildcard vmul.vx = {32'b100101_?_?????_?????_110_?????_1010111};
wildcard vmulh.vv = {32'b100111_?_?????_?????_010_?????_1010111};
wildcard vmulh.vx = {32'b100111_?_?????_?????_110_?????_1010111};
wildcard vmulhu.vv = {32'b100100_?_?????_?????_010_?????_1010111};
wildcard vmulhu.vx = {32'b100100_?_?????_?????_110_?????_1010111};
wildcard vmulhsu.vv = {32'b100110_?_?????_?????_010_?????_1010111};
wildcard vmulhsu.vx = {32'b100110_?_?????_?????_110_?????_1010111};
wildcard vdivu.vv = {32'b100000_?_?????_?????_010_?????_1010111};
wildcard vdivu.vx = {32'b100000_?_?????_?????_110_?????_1010111};
wildcard vdiv.vv = {32'b100001_?_?????_?????_010_?????_1010111};
wildcard vdiv.vx = {32'b100001_?_?????_?????_110_?????_1010111};
wildcard vremu.vv = {32'b100010_?_?????_?????_010_?????_1010111};
wildcard vremu.vx = {32'b100010_?_?????_?????_110_?????_1010111};
wildcard vrem.vv = {32'b100011_?_?????_?????_010_?????_1010111};
wildcard vrem.vx = {32'b100011_?_?????_?????_110_?????_1010111};
wildcard vwmul.vv = {32'b111011_?_?????_?????_010_?????_1010111};
wildcard vwmul.vx = {32'b111011_?_?????_?????_110_?????_1010111};
wildcard vwmulu.vv = {32'b111000_?_?????_?????_010_?????_1010111};
wildcard vwmulu.vx = {32'b111000_?_?????_?????_110_?????_1010111};
wildcard vwmulsu.vv = {32'b111010_?_?????_?????_010_?????_1010111};
wildcard vwmulsu.vx = {32'b111010_?_?????_?????_110_?????_1010111};
wildcard vmacc.vv = {32'b101101_?_?????_?????_010_?????_1010111};
wildcard vmacc.vx = {32'b101101_?_?????_?????_110_?????_1010111};
wildcard vnmsac.vv = {32'b101111_?_?????_?????_010_?????_1010111};
wildcard vnmsac.vx = {32'b101111_?_?????_?????_110_?????_1010111};
wildcard vmadd.vv = {32'b101001_?_?????_?????_010_?????_1010111};
wildcard vmadd.vx = {32'b101001_?_?????_?????_110_?????_1010111};
wildcard vnmsub.vv = {32'b101011_?_?????_?????_010_?????_1010111};
wildcard vnmsub.vx = {32'b101011_?_?????_?????_110_?????_1010111};
wildcard vwmaccu.vv = {32'b111100_?_?????_?????_010_?????_1010111};
wildcard vwmaccu.vx = {32'b111100_?_?????_?????_110_?????_1010111};
wildcard vwmacc.vv = {32'b111101_?_?????_?????_010_?????_1010111};
wildcard vwmacc.vx = {32'b111101_?_?????_?????_110_?????_1010111};
wildcard vwmaccsu.vv = {32'b111111_?_?????_?????_010_?????_1010111};
wildcard vwmaccsu.vx = {32'b111111_?_?????_?????_110_?????_1010111};
wildcard vwmaccus.vx = {32'b111110_?_?????_?????_110_?????_1010111};
wildcard vmerge.vvm = {32'b010111_0_?????_?????_000_?????_1010111};
wildcard vmerge.vxm = {32'b010111_0_?????_?????_100_?????_1010111};
wildcard vmerge.vim = {32'b010111_0_?????_?????_011_?????_1010111};
wildcard vmv.v.v = {32'b010111_1_00000_?????_000_?????_1010111};
wildcard vmv.v.x = {32'b010111_1_00000_?????_100_?????_1010111};
wildcard vmv.v.i = {32'b010111_1_00000_?????_011_?????_1010111};
wildcard vsaddu.vv = {32'b100000_?_?????_?????_000_?????_1010111};
wildcard vsaddu.vx = {32'b100000_?_?????_?????_100_?????_1010111};
wildcard vsaddu.vi = {32'b100000_?_?????_?????_011_?????_1010111};
wildcard vsadd.vv = {32'b100001_?_?????_?????_000_?????_1010111};
wildcard vsadd.vx = {32'b100001_?_?????_?????_100_?????_1010111};
wildcard vsadd.vi = {32'b100001_?_?????_?????_011_?????_1010111};
wildcard vssubu.vv = {32'b100010_?_?????_?????_000_?????_1010111};
wildcard vssubu.vx = {32'b100010_?_?????_?????_100_?????_1010111};
wildcard vssub.vv = {32'b100011_?_?????_?????_000_?????_1010111};
wildcard vssub.vx = {32'b100011_?_?????_?????_100_?????_1010111};
wildcard vaaddu.vv = {32'b001000_?_?????_?????_010_?????_1010111};
wildcard vaaddu.vx = {32'b001000_?_?????_?????_110_?????_1010111};
wildcard vaadd.vv = {32'b001001_?_?????_?????_010_?????_1010111};
wildcard vaadd.vx = {32'b001001_?_?????_?????_110_?????_1010111};
wildcard vasubu.vv = {32'b001010_?_?????_?????_010_?????_1010111};
wildcard vasubu.vx = {32'b001010_?_?????_?????_110_?????_1010111};
wildcard vasub.vv = {32'b001011_?_?????_?????_010_?????_1010111};
wildcard vasub.vx = {32'b001011_?_?????_?????_110_?????_1010111};
wildcard vsmul.vv = {32'b100111_?_?????_?????_000_?????_1010111};
wildcard vsmul.vx = {32'b100111_?_?????_?????_100_?????_1010111};
wildcard vssrl.vv = {32'b101010_?_?????_?????_000_?????_1010111};
wildcard vssrl.vx = {32'b101010_?_?????_?????_100_?????_1010111};
wildcard vssrl.vi = {32'b101010_?_?????_?????_011_?????_1010111};
wildcard vssra.vv = {32'b101011_?_?????_?????_000_?????_1010111};
wildcard vssra.vx = {32'b101011_?_?????_?????_100_?????_1010111};
wildcard vssra.vi = {32'b101011_?_?????_?????_011_?????_1010111};
wildcard vnclipu.wv = {32'b101110_?_?????_?????_000_?????_1010111};
wildcard vnclipu.wx = {32'b101110_?_?????_?????_100_?????_1010111};
wildcard vnclipu.wi = {32'b101110_?_?????_?????_011_?????_1010111};
wildcard vnclip.wv = {32'b101111_?_?????_?????_000_?????_1010111};
wildcard vnclip.wx = {32'b101111_?_?????_?????_100_?????_1010111};
wildcard vnclip.wi = {32'b101111_?_?????_?????_011_?????_1010111};
wildcard vfadd.vv = {32'b000000_?_?????_?????_001_?????_1010111};
wildcard vfadd.vf = {32'b000000_?_?????_?????_101_?????_1010111};
wildcard vfsub.vv = {32'b000010_?_?????_?????_001_?????_1010111};
wildcard vfsub.vf = {32'b000010_?_?????_?????_101_?????_1010111};
wildcard vfrsub.vf = {32'b100111_?_?????_?????_101_?????_1010111};
wildcard vfwadd.vv = {32'b110000_?_?????_?????_001_?????_1010111};
wildcard vfwadd.vf = {32'b110000_?_?????_?????_101_?????_1010111};
wildcard vfwsub.vv = {32'b110010_?_?????_?????_001_?????_1010111};
wildcard vfwsub.vf = {32'b110010_?_?????_?????_101_?????_1010111};
wildcard vfwadd.wv = {32'b110100_?_?????_?????_001_?????_1010111};
wildcard vfwadd.wf = {32'b110100_?_?????_?????_101_?????_1010111};
wildcard vfwsub.wv = {32'b110110_?_?????_?????_001_?????_1010111};
wildcard vfwsub.wf = {32'b110110_?_?????_?????_101_?????_1010111};
wildcard vfmul.vv = {32'b100100_?_?????_?????_001_?????_1010111};
wildcard vfmul.vf = {32'b100100_?_?????_?????_101_?????_1010111};
wildcard vfdiv.vv = {32'b100000_?_?????_?????_001_?????_1010111};
wildcard vfdiv.vf = {32'b100000_?_?????_?????_101_?????_1010111};
wildcard vfrdiv.vf = {32'b100001_?_?????_?????_101_?????_1010111};
wildcard vfwmul.vv = {32'b111000_?_?????_?????_001_?????_1010111};
wildcard vfwmul.vf = {32'b111000_?_?????_?????_101_?????_1010111};
wildcard vfmacc.vv = {32'b101100_?_?????_?????_001_?????_1010111};
wildcard vfmacc.vf = {32'b101100_?_?????_?????_101_?????_1010111};
wildcard vfnmacc.vv = {32'b101101_?_?????_?????_001_?????_1010111};
wildcard vfnmacc.vf = {32'b101101_?_?????_?????_101_?????_1010111};
wildcard vfmsac.vv = {32'b101110_?_?????_?????_001_?????_1010111};
wildcard vfmsac.vf = {32'b101110_?_?????_?????_101_?????_1010111};
wildcard vfnmsac.vv = {32'b101111_?_?????_?????_001_?????_1010111};
wildcard vfnmsac.vf = {32'b101111_?_?????_?????_101_?????_1010111};
wildcard vfmadd.vv = {32'b101000_?_?????_?????_001_?????_1010111};
wildcard vfmadd.vf = {32'b101000_?_?????_?????_101_?????_1010111};
wildcard vfnmadd.vv = {32'b101001_?_?????_?????_001_?????_1010111};
wildcard vfnmadd.vf = {32'b101001_?_?????_?????_101_?????_1010111};
wildcard vfmsub.vv = {32'b101010_?_?????_?????_001_?????_1010111};
wildcard vfmsub.vf = {32'b101010_?_?????_?????_101_?????_1010111};
wildcard vfnmsub.vv = {32'b101011_?_?????_?????_001_?????_1010111};
wildcard vfnmsub.vf = {32'b101011_?_?????_?????_101_?????_1010111};
wildcard vfwmacc.vv = {32'b111100_?_?????_?????_001_?????_1010111};
wildcard vfwmacc.vf = {32'b111100_?_?????_?????_101_?????_1010111};
wildcard vfwnmacc.vv = {32'b111101_?_?????_?????_001_?????_1010111};
wildcard vfwnmacc.vf = {32'b111101_?_?????_?????_101_?????_1010111};
wildcard vfwmsac.vv = {32'b111110_?_?????_?????_001_?????_1010111};
wildcard vfwmsac.vf = {32'b111110_?_?????_?????_101_?????_1010111};
wildcard vfwnmsac.vv = {32'b111111_?_?????_?????_001_?????_1010111};
wildcard vfwnmsac.vf = {32'b111111_?_?????_?????_101_?????_1010111};
wildcard vfsqrt.v = {32'b010011_?_?????_00000_001_?????_1010111};
wildcard vfrsqrt7.v = {32'b010011_?_?????_00100_001_?????_1010111};
wildcard vfrec7.v = {32'b010011_?_?????_00101_001_?????_1010111};
wildcard vfmin.vv = {32'b000100_?_?????_?????_001_?????_1010111};
wildcard vfmin.vf = {32'b000100_?_?????_?????_101_?????_1010111};
wildcard vfmax.vv = {32'b000110_?_?????_?????_001_?????_1010111};
wildcard vfmax.vf = {32'b000110_?_?????_?????_101_?????_1010111};
wildcard vfsgnj.vv = {32'b001000_?_?????_?????_001_?????_1010111};
wildcard vfsgnj.vf = {32'b001000_?_?????_?????_101_?????_1010111};
wildcard vfsgnjn.vv = {32'b001001_?_?????_?????_001_?????_1010111};
wildcard vfsgnjn.vf = {32'b001001_?_?????_?????_101_?????_1010111};
wildcard vfsgnjx.vv = {32'b001010_?_?????_?????_001_?????_1010111};
wildcard vfsgnjx.vf = {32'b001010_?_?????_?????_101_?????_1010111};
wildcard vmfeq.vv = {32'b011000_?_?????_?????_001_?????_1010111};
wildcard vmfeq.vf = {32'b011000_?_?????_?????_101_?????_1010111};
wildcard vmfne.vv = {32'b011100_?_?????_?????_001_?????_1010111};
wildcard vmfne.vf = {32'b011100_?_?????_?????_101_?????_1010111};
wildcard vmflt.vv = {32'b011011_?_?????_?????_001_?????_1010111};
wildcard vmflt.vf = {32'b011011_?_?????_?????_101_?????_1010111};
wildcard vmfle.vv = {32'b011001_?_?????_?????_001_?????_1010111};
wildcard vmfle.vf = {32'b011001_?_?????_?????_101_?????_1010111};
wildcard vmfgt.vf = {32'b011101_?_?????_?????_101_?????_1010111};
wildcard vmfge.vf = {32'b011111_?_?????_?????_101_?????_1010111};
wildcard vfclass.v = {32'b010011_?_?????_10000_001_?????_1010111};
wildcard vfmerge.vfm = {32'b010111_?_?????_?????_101_?????_1010111};
wildcard vfmv.v.f = {32'b010111_?_?????_?????_101_?????_1010111};
wildcard vfcvt.xu.f.v = {32'b010010_?_?????_00000_001_?????_1010111};
wildcard vfcvt.x.f.v = {32'b010010_?_?????_00001_001_?????_1010111};
wildcard vfcvt.rtz.xu.f.v = {32'b010010_?_?????_00110_001_?????_1010111};
wildcard vfcvt.rtz.x.f.v = {32'b010010_?_?????_00111_001_?????_1010111};
wildcard vfcvt.f.xu.v = {32'b010010_?_?????_00010_001_?????_1010111};
wildcard vfcvt.f.x.v = {32'b010010_?_?????_00011_001_?????_1010111};
wildcard vfwcvt.xu.f.v = {32'b010010_?_?????_01000_001_?????_1010111};
wildcard vfwcvt.x.f.v = {32'b010010_?_?????_01001_001_?????_1010111};
wildcard vfwcvt.rtz.xu.f.v = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfwcvt.rtz.x.f.v = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfwcvt.f.xu.v = {32'b010010_?_?????_01010_001_?????_1010111};
wildcard vfwcvt.f.x.v = {32'b010010_?_?????_01011_001_?????_1010111};
wildcard vfwcvt.f.f.v = {32'b010010_?_?????_01100_001_?????_1010111};
wildcard vfncvt.xu.f.w = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfncvt.x.f.w = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfncvt.rtz.xu.f.w = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfncvt.rtz.x.f.w = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfncvt.f.xu.w = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfncvt.f.x.w = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfncvt.f.f.w = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vfncvt.rod.f.f.w = {32'b010010_?_?????_?????_001_?????_1010111};
wildcard vredsum.vs = {32'b000000_?_?????_?????_010_?????_1010111};
wildcard vredmaxu.vs = {32'b000110_?_?????_?????_010_?????_1010111};
wildcard vredmax.vs = {32'b000111_?_?????_?????_010_?????_1010111};
wildcard vredminu.vs = {32'b000100_?_?????_?????_010_?????_1010111};
wildcard vredmin.vs = {32'b000101_?_?????_?????_010_?????_1010111};
wildcard vredand.vs = {32'b000001_?_?????_?????_010_?????_1010111};
wildcard vredor.vs = {32'b000011_?_?????_?????_010_?????_1010111};
wildcard vredxor.vs = {32'b000011_?_?????_?????_010_?????_1010111};
wildcard vwredsumu.vs = {32'b110000_?_?????_?????_000_?????_1010111};
wildcard vwredsum.vs = {32'b110001_?_?????_?????_000_?????_1010111};
wildcard vfredosum.vs = {32'b000011_?_?????_?????_001_?????_1010111};
wildcard vfredusum.vs = {32'b000001_?_?????_?????_001_?????_1010111};
wildcard vfredmax.vs = {32'b000111_?_?????_?????_001_?????_1010111};
wildcard vfredmin.vs = {32'b000101_?_?????_?????_001_?????_1010111};
wildcard vfwredosum.vs = {32'b110011_?_?????_?????_001_?????_1010111};
wildcard vfwredusum.vs = {32'b110001_?_?????_?????_001_?????_1010111};
wildcard vmand.mm = {32'b011001_?_?????_?????_010_?????_1010111};
wildcard vmnand.mm = {32'b011101_?_?????_?????_010_?????_1010111};
wildcard vmandn.mm = {32'b011000_?_?????_?????_010_?????_1010111};
wildcard vmxor.mm = {32'b011011_?_?????_?????_010_?????_1010111};
wildcard vmor.mm = {32'b011010_?_?????_?????_010_?????_1010111};
wildcard vmnor.mm = {32'b011110_?_?????_?????_010_?????_1010111};
wildcard vmorn.mm = {32'b011100_?_?????_?????_010_?????_1010111};
wildcard vmxnor.mm = {32'b011111_?_?????_?????_010_?????_1010111};
wildcard vcpop.m = {32'b010000_?_?????_10000_010_?????_1010111};
wildcard vfirst.m = {32'b010000_?_?????_10001_010_?????_1010111};
wildcard vmsbf.m = {32'b010100_?_?????_00001_010_?????_1010111};
wildcard vmsif.m = {32'b010100_?_?????_00011_010_?????_1010111};
wildcard vmsof.m = {32'b010100_?_?????_00010_010_?????_1010111};
wildcard viota.m = {32'b010100_?_?????_10000_010_?????_1010111};
wildcard vid.v = {32'b010100_?_?????_10001_010_?????_1010111};
wildcard vmv.x.s = {32'b010000_?_?????_000000_010_?????_1010111};
wildcard vmv.s.x = {32'b010000_?_00000_?????_110_?????_1010111};
wildcard vfmv.f.s = {32'b010000_?_?????_00000_001_?????_1010111};
wildcard vfmv.s.f = {32'b010000_?_?????_?????_101_?????_1010111};
wildcard vslideup.vx = {32'b001110_?_?????_?????_100_?????_1010111};
wildcard vslideup.vi = {32'b001110_?_?????_?????_011_?????_1010111};
wildcard vslidedown.vx = {32'b001111_?_?????_?????_100_?????_1010111};
wildcard vslidedown.vi = {32'b001111_?_?????_?????_011_?????_1010111};
wildcard vslide1up.vx = {32'b001110_?_?????_?????_110_?????_1010111};
wildcard vfslide1up.vf = {32'b001110_?_?????_?????_101_?????_1010111};
wildcard vslide1down.vx = {32'b001111_?_?????_?????_110_?????_1010111};
wildcard vfslide1down.vf = {32'b001111_?_?????_?????_101_?????_1010111};
wildcard vrgather.vv = {32'b001100_?_?????_?????_000_?????_1010111};
wildcard vrgatherei16.vv = {32'b001110_?_?????_?????_000_?????_1010111};
wildcard vrgather.vx = {32'b001100_?_?????_?????_100_?????_1010111};
wildcard vrgather.vi = {32'b001100_?_?????_?????_011_?????_1010111};
wildcard vcompress.vm = {32'b010111_?_?????_?????_010_?????_1010111};
wildcard vmv1r.v = {32'b100111_1_?????_??000_011_?????_1010111};
wildcard vmv2r.v = {32'b100111_1_?????_??001_011_?????_1010111};
wildcard vmv4r.v = {32'b100111_1_?????_??011_011_?????_1010111};
wildcard vmv8r.v = {32'b100111_1_?????_??110_011_?????_1010111};
