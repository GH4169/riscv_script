wildcard vadd_OPIVV = {32'b000000_?_?????_?????_000_?????_1010111};
wildcard vadd_OPIVX = {32'b000000_?_?????_?????_100_?????_1010111};
wildcard vadd_OPIVI = {32'b000000_?_?????_?????_011_?????_1010111};
wildcard vsub_OPIVV = {32'b000010_?_?????_?????_000_?????_1010111};
wildcard vsub_OPIVX = {32'b000010_?_?????_?????_100_?????_1010111};
wildcard vrsub_OPIVX = {32'b000011_?_?????_?????_100_?????_1010111};
wildcard vrsub_OPIVI = {32'b000011_?_?????_?????_011_?????_1010111};
wildcard vminu_OPIVV = {32'b000100_?_?????_?????_000_?????_1010111};
wildcard vminu_OPIVX = {32'b000100_?_?????_?????_100_?????_1010111};
wildcard vmin_OPIVV = {32'b000101_?_?????_?????_000_?????_1010111};
wildcard vmin_OPIVX = {32'b000101_?_?????_?????_100_?????_1010111};
wildcard vmaxu_OPIVV = {32'b000110_?_?????_?????_000_?????_1010111};
wildcard vmaxu_OPIVX = {32'b000110_?_?????_?????_100_?????_1010111};
wildcard vmax_OPIVV = {32'b000111_?_?????_?????_000_?????_1010111};
wildcard vmax_OPIVX = {32'b000111_?_?????_?????_100_?????_1010111};
wildcard vand_OPIVV = {32'b001001_?_?????_?????_000_?????_1010111};
wildcard vand_OPIVX = {32'b001001_?_?????_?????_100_?????_1010111};
wildcard vand_OPIVI = {32'b001001_?_?????_?????_011_?????_1010111};
wildcard vor_OPIVV = {32'b001010_?_?????_?????_000_?????_1010111};
wildcard vor_OPIVX = {32'b001010_?_?????_?????_100_?????_1010111};
wildcard vor_OPIVI = {32'b001010_?_?????_?????_011_?????_1010111};
wildcard vxor_OPIVV = {32'b001011_?_?????_?????_000_?????_1010111};
wildcard vxor_OPIVX = {32'b001011_?_?????_?????_100_?????_1010111};
wildcard vxor_OPIVI = {32'b001011_?_?????_?????_011_?????_1010111};
wildcard vrgather_OPIVV = {32'b001100_?_?????_?????_000_?????_1010111};
wildcard vrgather_OPIVX = {32'b001100_?_?????_?????_100_?????_1010111};
wildcard vrgather_OPIVI = {32'b001100_?_?????_?????_011_?????_1010111};
wildcard vslideup_OPIVX = {32'b001110_?_?????_?????_100_?????_1010111};
wildcard vslideup_OPIVI = {32'b001110_?_?????_?????_011_?????_1010111};
wildcard vrgatherei16_OPIVV = {32'b001110_?_?????_?????_000_?????_1010111};
wildcard vslidedown_OPIVX = {32'b001111_?_?????_?????_100_?????_1010111};
wildcard vslidedown_OPIVI = {32'b001111_?_?????_?????_011_?????_1010111};
wildcard vadc_OPIVV = {32'b010000_?_?????_?????_000_?????_1010111};
wildcard vadc_OPIVX = {32'b010000_?_?????_?????_100_?????_1010111};
wildcard vadc_OPIVI = {32'b010000_?_?????_?????_011_?????_1010111};
wildcard vmadc_OPIVV = {32'b010001_?_?????_?????_000_?????_1010111};
wildcard vmadc_OPIVX = {32'b010001_?_?????_?????_100_?????_1010111};
wildcard vmadc_OPIVI = {32'b010001_?_?????_?????_011_?????_1010111};
wildcard vsbc_OPIVV = {32'b010010_?_?????_?????_000_?????_1010111};
wildcard vsbc_OPIVX = {32'b010010_?_?????_?????_100_?????_1010111};
wildcard vmsbc_OPIVV = {32'b010011_?_?????_?????_000_?????_1010111};
wildcard vmsbc_OPIVX = {32'b010011_?_?????_?????_100_?????_1010111};
wildcard vmerge/vmv_OPIVV = {32'b010111_?_?????_?????_000_?????_1010111};
wildcard vmerge/vmv_OPIVX = {32'b010111_?_?????_?????_100_?????_1010111};
wildcard vmerge/vmv_OPIVI = {32'b010111_?_?????_?????_011_?????_1010111};
wildcard vmseq_OPIVV = {32'b011000_?_?????_?????_000_?????_1010111};
wildcard vmseq_OPIVX = {32'b011000_?_?????_?????_100_?????_1010111};
wildcard vmseq_OPIVI = {32'b011000_?_?????_?????_011_?????_1010111};
wildcard vmsne_OPIVV = {32'b011001_?_?????_?????_000_?????_1010111};
wildcard vmsne_OPIVX = {32'b011001_?_?????_?????_100_?????_1010111};
wildcard vmsne_OPIVI = {32'b011001_?_?????_?????_011_?????_1010111};
wildcard vmsltu_OPIVV = {32'b011010_?_?????_?????_000_?????_1010111};
wildcard vmsltu_OPIVX = {32'b011010_?_?????_?????_100_?????_1010111};
wildcard vmslt_OPIVV = {32'b011011_?_?????_?????_000_?????_1010111};
wildcard vmslt_OPIVX = {32'b011011_?_?????_?????_100_?????_1010111};
wildcard vmsleu_OPIVV = {32'b011100_?_?????_?????_000_?????_1010111};
wildcard vmsleu_OPIVX = {32'b011100_?_?????_?????_100_?????_1010111};
wildcard vmsleu_OPIVI = {32'b011100_?_?????_?????_011_?????_1010111};
wildcard vmsle_OPIVV = {32'b011101_?_?????_?????_000_?????_1010111};
wildcard vmsle_OPIVX = {32'b011101_?_?????_?????_100_?????_1010111};
wildcard vmsle_OPIVI = {32'b011101_?_?????_?????_011_?????_1010111};
wildcard vmsgtu_OPIVX = {32'b011110_?_?????_?????_100_?????_1010111};
wildcard vmsgtu_OPIVI = {32'b011110_?_?????_?????_011_?????_1010111};
wildcard vmsgt_OPIVX = {32'b011111_?_?????_?????_100_?????_1010111};
wildcard vmsgt_OPIVI = {32'b011111_?_?????_?????_011_?????_1010111};
wildcard vsaddu_OPIVV = {32'b100000_?_?????_?????_000_?????_1010111};
wildcard vsaddu_OPIVX = {32'b100000_?_?????_?????_100_?????_1010111};
wildcard vsaddu_OPIVI = {32'b100000_?_?????_?????_011_?????_1010111};
wildcard vsadd_OPIVV = {32'b100001_?_?????_?????_000_?????_1010111};
wildcard vsadd_OPIVX = {32'b100001_?_?????_?????_100_?????_1010111};
wildcard vsadd_OPIVI = {32'b100001_?_?????_?????_011_?????_1010111};
wildcard vssubu_OPIVV = {32'b100010_?_?????_?????_000_?????_1010111};
wildcard vssubu_OPIVX = {32'b100010_?_?????_?????_100_?????_1010111};
wildcard vssub_OPIVV = {32'b100011_?_?????_?????_000_?????_1010111};
wildcard vssub_OPIVX = {32'b100011_?_?????_?????_100_?????_1010111};
wildcard vsll_OPIVV = {32'b100101_?_?????_?????_000_?????_1010111};
wildcard vsll_OPIVX = {32'b100101_?_?????_?????_100_?????_1010111};
wildcard vsll_OPIVI = {32'b100101_?_?????_?????_011_?????_1010111};
wildcard vsmul_OPIVV = {32'b100111_?_?????_?????_000_?????_1010111};
wildcard vsmul_OPIVX = {32'b100111_?_?????_?????_100_?????_1010111};
wildcard vmv<nr>r_OPIVI = {32'b100111_?_?????_?????_011_?????_1010111};
wildcard vsrl_OPIVV = {32'b101000_?_?????_?????_000_?????_1010111};
wildcard vsrl_OPIVX = {32'b101000_?_?????_?????_100_?????_1010111};
wildcard vsrl_OPIVI = {32'b101000_?_?????_?????_011_?????_1010111};
wildcard vsra_OPIVV = {32'b101001_?_?????_?????_000_?????_1010111};
wildcard vsra_OPIVX = {32'b101001_?_?????_?????_100_?????_1010111};
wildcard vsra_OPIVI = {32'b101001_?_?????_?????_011_?????_1010111};
wildcard vssrl_OPIVV = {32'b101010_?_?????_?????_000_?????_1010111};
wildcard vssrl_OPIVX = {32'b101010_?_?????_?????_100_?????_1010111};
wildcard vssrl_OPIVI = {32'b101010_?_?????_?????_011_?????_1010111};
wildcard vssra_OPIVV = {32'b101011_?_?????_?????_000_?????_1010111};
wildcard vssra_OPIVX = {32'b101011_?_?????_?????_100_?????_1010111};
wildcard vssra_OPIVI = {32'b101011_?_?????_?????_011_?????_1010111};
wildcard vnsrl_OPIVV = {32'b101100_?_?????_?????_000_?????_1010111};
wildcard vnsrl_OPIVX = {32'b101100_?_?????_?????_100_?????_1010111};
wildcard vnsrl_OPIVI = {32'b101100_?_?????_?????_011_?????_1010111};
wildcard vnsra_OPIVV = {32'b101101_?_?????_?????_000_?????_1010111};
wildcard vnsra_OPIVX = {32'b101101_?_?????_?????_100_?????_1010111};
wildcard vnsra_OPIVI = {32'b101101_?_?????_?????_011_?????_1010111};
wildcard vnclipu_OPIVV = {32'b101110_?_?????_?????_000_?????_1010111};
wildcard vnclipu_OPIVX = {32'b101110_?_?????_?????_100_?????_1010111};
wildcard vnclipu_OPIVI = {32'b101110_?_?????_?????_011_?????_1010111};
wildcard vnclip_OPIVV = {32'b101111_?_?????_?????_000_?????_1010111};
wildcard vnclip_OPIVX = {32'b101111_?_?????_?????_100_?????_1010111};
wildcard vnclip_OPIVI = {32'b101111_?_?????_?????_011_?????_1010111};
wildcard vwredsumu_OPIVV = {32'b110000_?_?????_?????_000_?????_1010111};
wildcard vwredsum_OPIVV = {32'b110001_?_?????_?????_000_?????_1010111};
wildcard vredsum_OPMVV = {32'b000000_?_?????_?????_010_?????_1010111};
wildcard vredand_OPMVV = {32'b000001_?_?????_?????_010_?????_1010111};
wildcard vredor_OPMVV = {32'b000010_?_?????_?????_010_?????_1010111};
wildcard vredxor_OPMVV = {32'b000011_?_?????_?????_010_?????_1010111};
wildcard vredminu_OPMVV = {32'b000100_?_?????_?????_010_?????_1010111};
wildcard vredmin_OPMVV = {32'b000101_?_?????_?????_010_?????_1010111};
wildcard vredmaxu_OPMVV = {32'b000110_?_?????_?????_010_?????_1010111};
wildcard vredmax_OPMVV = {32'b000111_?_?????_?????_010_?????_1010111};
wildcard vaaddu_OPMVV = {32'b001000_?_?????_?????_010_?????_1010111};
wildcard vaaddu_OPMVX = {32'b001000_?_?????_?????_110_?????_1010111};
wildcard vaadd_OPMVV = {32'b001001_?_?????_?????_010_?????_1010111};
wildcard vaadd_OPMVX = {32'b001001_?_?????_?????_110_?????_1010111};
wildcard vasubu_OPMVV = {32'b001010_?_?????_?????_010_?????_1010111};
wildcard vasubu_OPMVX = {32'b001010_?_?????_?????_110_?????_1010111};
wildcard vasub_OPMVV = {32'b001011_?_?????_?????_010_?????_1010111};
wildcard vasub_OPMVX = {32'b001011_?_?????_?????_110_?????_1010111};
wildcard vslide1up_OPMVX = {32'b001110_?_?????_?????_110_?????_1010111};
wildcard vslide1down_OPMVX = {32'b001111_?_?????_?????_110_?????_1010111};
wildcard vcompress_OPMVV = {32'b010111_?_?????_?????_010_?????_1010111};
wildcard vmandn_OPMVV = {32'b011000_?_?????_?????_010_?????_1010111};
wildcard vmand_OPMVV = {32'b011001_?_?????_?????_010_?????_1010111};
wildcard vmor_OPMVV = {32'b011010_?_?????_?????_010_?????_1010111};
wildcard vmxor_OPMVV = {32'b011011_?_?????_?????_010_?????_1010111};
wildcard vmorn_OPMVV = {32'b011100_?_?????_?????_010_?????_1010111};
wildcard vmnand_OPMVV = {32'b011101_?_?????_?????_010_?????_1010111};
wildcard vmnor_OPMVV = {32'b011110_?_?????_?????_010_?????_1010111};
wildcard vmxnor_OPMVV = {32'b011111_?_?????_?????_010_?????_1010111};
wildcard vdivu_OPMVV = {32'b100000_?_?????_?????_010_?????_1010111};
wildcard vdivu_OPMVX = {32'b100000_?_?????_?????_110_?????_1010111};
wildcard vdiv_OPMVV = {32'b100001_?_?????_?????_010_?????_1010111};
wildcard vdiv_OPMVX = {32'b100001_?_?????_?????_110_?????_1010111};
wildcard vremu_OPMVV = {32'b100010_?_?????_?????_010_?????_1010111};
wildcard vremu_OPMVX = {32'b100010_?_?????_?????_110_?????_1010111};
wildcard vrem_OPMVV = {32'b100011_?_?????_?????_010_?????_1010111};
wildcard vrem_OPMVX = {32'b100011_?_?????_?????_110_?????_1010111};
wildcard vmulhu_OPMVV = {32'b100100_?_?????_?????_010_?????_1010111};
wildcard vmulhu_OPMVX = {32'b100100_?_?????_?????_110_?????_1010111};
wildcard vmul_OPMVV = {32'b100101_?_?????_?????_010_?????_1010111};
wildcard vmul_OPMVX = {32'b100101_?_?????_?????_110_?????_1010111};
wildcard vmulhsu_OPMVV = {32'b100110_?_?????_?????_010_?????_1010111};
wildcard vmulhsu_OPMVX = {32'b100110_?_?????_?????_110_?????_1010111};
wildcard vmulh_OPMVV = {32'b100111_?_?????_?????_010_?????_1010111};
wildcard vmulh_OPMVX = {32'b100111_?_?????_?????_110_?????_1010111};
wildcard vmadd_OPMVV = {32'b101001_?_?????_?????_010_?????_1010111};
wildcard vmadd_OPMVX = {32'b101001_?_?????_?????_110_?????_1010111};
wildcard vnmsub_OPMVV = {32'b101011_?_?????_?????_010_?????_1010111};
wildcard vnmsub_OPMVX = {32'b101011_?_?????_?????_110_?????_1010111};
wildcard vmacc_OPMVV = {32'b101101_?_?????_?????_010_?????_1010111};
wildcard vmacc_OPMVX = {32'b101101_?_?????_?????_110_?????_1010111};
wildcard vnmsac_OPMVV = {32'b101111_?_?????_?????_010_?????_1010111};
wildcard vnmsac_OPMVX = {32'b101111_?_?????_?????_110_?????_1010111};
wildcard vwaddu_OPMVV = {32'b110000_?_?????_?????_010_?????_1010111};
wildcard vwaddu_OPMVX = {32'b110000_?_?????_?????_110_?????_1010111};
wildcard vwadd_OPMVV = {32'b110001_?_?????_?????_010_?????_1010111};
wildcard vwadd_OPMVX = {32'b110001_?_?????_?????_110_?????_1010111};
wildcard vwsubu_OPMVV = {32'b110010_?_?????_?????_010_?????_1010111};
wildcard vwsubu_OPMVX = {32'b110010_?_?????_?????_110_?????_1010111};
wildcard vwsub_OPMVV = {32'b110011_?_?????_?????_010_?????_1010111};
wildcard vwsub_OPMVX = {32'b110011_?_?????_?????_110_?????_1010111};
wildcard vwaddu.w_OPMVV = {32'b110100_?_?????_?????_010_?????_1010111};
wildcard vwaddu.w_OPMVX = {32'b110100_?_?????_?????_110_?????_1010111};
wildcard vwadd.w_OPMVV = {32'b110101_?_?????_?????_010_?????_1010111};
wildcard vwadd.w_OPMVX = {32'b110101_?_?????_?????_110_?????_1010111};
wildcard vwsubu.w_OPMVV = {32'b110110_?_?????_?????_010_?????_1010111};
wildcard vwsubu.w_OPMVX = {32'b110110_?_?????_?????_110_?????_1010111};
wildcard vwsub.w_OPMVV = {32'b110111_?_?????_?????_010_?????_1010111};
wildcard vwsub.w_OPMVX = {32'b110111_?_?????_?????_110_?????_1010111};
wildcard vwmulu_OPMVV = {32'b111000_?_?????_?????_010_?????_1010111};
wildcard vwmulu_OPMVX = {32'b111000_?_?????_?????_110_?????_1010111};
wildcard vwmulsu_OPMVV = {32'b111010_?_?????_?????_010_?????_1010111};
wildcard vwmulsu_OPMVX = {32'b111010_?_?????_?????_110_?????_1010111};
wildcard vwmul_OPMVV = {32'b111011_?_?????_?????_010_?????_1010111};
wildcard vwmul_OPMVX = {32'b111011_?_?????_?????_110_?????_1010111};
wildcard vwmaccu_OPMVV = {32'b111100_?_?????_?????_010_?????_1010111};
wildcard vwmaccu_OPMVX = {32'b111100_?_?????_?????_110_?????_1010111};
wildcard vwmacc_OPMVV = {32'b111101_?_?????_?????_010_?????_1010111};
wildcard vwmacc_OPMVX = {32'b111101_?_?????_?????_110_?????_1010111};
wildcard vwmaccus_OPMVX = {32'b111110_?_?????_?????_110_?????_1010111};
wildcard vwmaccsu_OPMVV = {32'b111111_?_?????_?????_010_?????_1010111};
wildcard vwmaccsu_OPMVX = {32'b111111_?_?????_?????_110_?????_1010111};
wildcard vfadd_OPFVV = {32'b000000_?_?????_?????_001_?????_1010111};
wildcard vfadd_OPFVF = {32'b000000_?_?????_?????_101_?????_1010111};
wildcard vfredusum_OPFVV = {32'b000001_?_?????_?????_001_?????_1010111};
wildcard vfsub_OPFVV = {32'b000010_?_?????_?????_001_?????_1010111};
wildcard vfsub_OPFVF = {32'b000010_?_?????_?????_101_?????_1010111};
wildcard vfredosum_OPFVV = {32'b000011_?_?????_?????_001_?????_1010111};
wildcard vfmin_OPFVV = {32'b000100_?_?????_?????_001_?????_1010111};
wildcard vfmin_OPFVF = {32'b000100_?_?????_?????_101_?????_1010111};
wildcard vfredmin_OPFVV = {32'b000101_?_?????_?????_001_?????_1010111};
wildcard vfmax_OPFVV = {32'b000110_?_?????_?????_001_?????_1010111};
wildcard vfmax_OPFVF = {32'b000110_?_?????_?????_101_?????_1010111};
wildcard vfredmax_OPFVV = {32'b000111_?_?????_?????_001_?????_1010111};
wildcard vfsgnj_OPFVV = {32'b001000_?_?????_?????_001_?????_1010111};
wildcard vfsgnj_OPFVF = {32'b001000_?_?????_?????_101_?????_1010111};
wildcard vfsgnjn_OPFVV = {32'b001001_?_?????_?????_001_?????_1010111};
wildcard vfsgnjn_OPFVF = {32'b001001_?_?????_?????_101_?????_1010111};
wildcard vfsgnjx_OPFVV = {32'b001010_?_?????_?????_001_?????_1010111};
wildcard vfsgnjx_OPFVF = {32'b001010_?_?????_?????_101_?????_1010111};
wildcard vfslide1up_OPFVF = {32'b001110_?_?????_?????_101_?????_1010111};
wildcard vfslide1down_OPFVF = {32'b001111_?_?????_?????_101_?????_1010111};
wildcard vfmerge/vfmv_OPFVF = {32'b010111_?_?????_?????_101_?????_1010111};
wildcard vmfeq_OPFVV = {32'b011000_?_?????_?????_001_?????_1010111};
wildcard vmfeq_OPFVF = {32'b011000_?_?????_?????_101_?????_1010111};
wildcard vmfle_OPFVV = {32'b011001_?_?????_?????_001_?????_1010111};
wildcard vmfle_OPFVF = {32'b011001_?_?????_?????_101_?????_1010111};
wildcard vmflt_OPFVV = {32'b011011_?_?????_?????_001_?????_1010111};
wildcard vmflt_OPFVF = {32'b011011_?_?????_?????_101_?????_1010111};
wildcard vmfne_OPFVV = {32'b011100_?_?????_?????_001_?????_1010111};
wildcard vmfne_OPFVF = {32'b011100_?_?????_?????_101_?????_1010111};
wildcard vmfgt_OPFVF = {32'b011101_?_?????_?????_101_?????_1010111};
wildcard vmfge_OPFVF = {32'b011111_?_?????_?????_101_?????_1010111};
wildcard vfdiv_OPFVV = {32'b100000_?_?????_?????_001_?????_1010111};
wildcard vfdiv_OPFVF = {32'b100000_?_?????_?????_101_?????_1010111};
wildcard vfrdiv_OPFVF = {32'b100001_?_?????_?????_101_?????_1010111};
wildcard vfmul_OPFVV = {32'b100100_?_?????_?????_001_?????_1010111};
wildcard vfmul_OPFVF = {32'b100100_?_?????_?????_101_?????_1010111};
wildcard vfrsub_OPFVF = {32'b100111_?_?????_?????_101_?????_1010111};
wildcard vfmadd_OPFVV = {32'b101000_?_?????_?????_001_?????_1010111};
wildcard vfmadd_OPFVF = {32'b101000_?_?????_?????_101_?????_1010111};
wildcard vfnmadd_OPFVV = {32'b101001_?_?????_?????_001_?????_1010111};
wildcard vfnmadd_OPFVF = {32'b101001_?_?????_?????_101_?????_1010111};
wildcard vfmsub_OPFVV = {32'b101010_?_?????_?????_001_?????_1010111};
wildcard vfmsub_OPFVF = {32'b101010_?_?????_?????_101_?????_1010111};
wildcard vfnmsub_OPFVV = {32'b101011_?_?????_?????_001_?????_1010111};
wildcard vfnmsub_OPFVF = {32'b101011_?_?????_?????_101_?????_1010111};
wildcard vfmacc_OPFVV = {32'b101100_?_?????_?????_001_?????_1010111};
wildcard vfmacc_OPFVF = {32'b101100_?_?????_?????_101_?????_1010111};
wildcard vfnmacc_OPFVV = {32'b101101_?_?????_?????_001_?????_1010111};
wildcard vfnmacc_OPFVF = {32'b101101_?_?????_?????_101_?????_1010111};
wildcard vfmsac_OPFVV = {32'b101110_?_?????_?????_001_?????_1010111};
wildcard vfmsac_OPFVF = {32'b101110_?_?????_?????_101_?????_1010111};
wildcard vfnmsac_OPFVV = {32'b101111_?_?????_?????_001_?????_1010111};
wildcard vfnmsac_OPFVF = {32'b101111_?_?????_?????_101_?????_1010111};
wildcard vfwadd_OPFVV = {32'b110000_?_?????_?????_001_?????_1010111};
wildcard vfwadd_OPFVF = {32'b110000_?_?????_?????_101_?????_1010111};
wildcard vfwredusum_OPFVV = {32'b110001_?_?????_?????_001_?????_1010111};
wildcard vfwsub_OPFVV = {32'b110010_?_?????_?????_001_?????_1010111};
wildcard vfwsub_OPFVF = {32'b110010_?_?????_?????_101_?????_1010111};
wildcard vfwredosum_OPFVV = {32'b110011_?_?????_?????_001_?????_1010111};
wildcard vfwadd.w_OPFVV = {32'b110100_?_?????_?????_001_?????_1010111};
wildcard vfwadd.w_OPFVF = {32'b110100_?_?????_?????_101_?????_1010111};
wildcard vfwsub.w_OPFVV = {32'b110110_?_?????_?????_001_?????_1010111};
wildcard vfwsub.w_OPFVF = {32'b110110_?_?????_?????_101_?????_1010111};
wildcard vfwmul_OPFVV = {32'b111000_?_?????_?????_001_?????_1010111};
wildcard vfwmul_OPFVF = {32'b111000_?_?????_?????_101_?????_1010111};
wildcard vfwmacc_OPFVV = {32'b111100_?_?????_?????_001_?????_1010111};
wildcard vfwmacc_OPFVF = {32'b111100_?_?????_?????_101_?????_1010111};
wildcard vfwnmacc_OPFVV = {32'b111101_?_?????_?????_001_?????_1010111};
wildcard vfwnmacc_OPFVF = {32'b111101_?_?????_?????_101_?????_1010111};
wildcard vfwmsac_OPFVV = {32'b111110_?_?????_?????_001_?????_1010111};
wildcard vfwmsac_OPFVF = {32'b111110_?_?????_?????_101_?????_1010111};
wildcard vfwnmsac_OPFVV = {32'b111111_?_?????_?????_001_?????_1010111};
wildcard vfwnmsac_OPFVF = {32'b111111_?_?????_?????_101_?????_1010111};
wildcard VRXUNARY0_OPMVX_rs2_vmv.s.x = {32'b010000_?_00000_?????_110_?????_1010111};
wildcard VWXUNARY0_OPMVV_rs1_vmv.x.s = {32'b010000_?_?????_00000_010_?????_1010111};
wildcard VWXUNARY0_OPMVV_rs1_vcpop = {32'b010000_?_?????_10000_010_?????_1010111};
wildcard VWXUNARY0_OPMVV_rs1_vfirst = {32'b010000_?_?????_10001_010_?????_1010111};
wildcard VXUNARY0_OPMVV_rs1_vzext.vf8 = {32'b010010_?_?????_00010_010_?????_1010111};
wildcard VXUNARY0_OPMVV_rs1_vsext.vf8 = {32'b010010_?_?????_00011_010_?????_1010111};
wildcard VXUNARY0_OPMVV_rs1_vzext.vf4 = {32'b010010_?_?????_00100_010_?????_1010111};
wildcard VXUNARY0_OPMVV_rs1_vsext.vf4 = {32'b010010_?_?????_00101_010_?????_1010111};
wildcard VXUNARY0_OPMVV_rs1_vzext.vf2 = {32'b010010_?_?????_00110_010_?????_1010111};
wildcard VXUNARY0_OPMVV_rs1_vsext.vf2 = {32'b010010_?_?????_00111_010_?????_1010111};
wildcard VRFUNARY0_OPFVF_rs2_vfmv.s.f = {32'b010000_?_00000_?????_101_?????_1010111};
wildcard VWFUNARY0_OPFVV_rs1_vfmv.f.s = {32'b010000_?_?????_00000_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfcvt.xu.f.v = {32'b010010_?_?????_00000_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfcvt.x.f.v = {32'b010010_?_?????_00001_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfcvt.f.xu.v = {32'b010010_?_?????_00010_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfcvt.f.x.v = {32'b010010_?_?????_00011_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfcvt.rtz.xu.f.v = {32'b010010_?_?????_00110_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfcvt.rtz.x.f.v = {32'b010010_?_?????_00111_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfwcvt.xu.f.v = {32'b010010_?_?????_01000_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfwcvt.x.f.v = {32'b010010_?_?????_01001_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfwcvt.f.xu.v = {32'b010010_?_?????_01010_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfwcvt.f.x.v = {32'b010010_?_?????_01011_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfwcvt.f.f.v = {32'b010010_?_?????_01100_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfwcvt.rtz.xu.f.v = {32'b010010_?_?????_01110_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfwcvt.rtz.x.f.v = {32'b010010_?_?????_01111_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfncvt.xu.f.w = {32'b010010_?_?????_10000_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfncvt.x.f.w = {32'b010010_?_?????_10001_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfncvt.f.xu.w = {32'b010010_?_?????_10010_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfncvt.f.x.w = {32'b010010_?_?????_10011_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfncvt.f.f.w = {32'b010010_?_?????_10100_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfncvt.rod.f.f.w = {32'b010010_?_?????_10101_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfncvt.rtz.xu.f.w = {32'b010010_?_?????_10110_001_?????_1010111};
wildcard VFUNARY0_OPFVV_rs1_vfncvt.rtz.x.f.w = {32'b010010_?_?????_10111_001_?????_1010111};
wildcard VFUNARY1_OPFVV_rs1_vfsqrt.v = {32'b010011_?_?????_00000_001_?????_1010111};
wildcard VFUNARY1_OPFVV_rs1_vfrsqrt7.v = {32'b010011_?_?????_00100_001_?????_1010111};
wildcard VFUNARY1_OPFVV_rs1_vfrec7.v = {32'b010011_?_?????_00101_001_?????_1010111};
wildcard VFUNARY1_OPFVV_rs1_vfclass.v = {32'b010011_?_?????_10000_001_?????_1010111};
wildcard VMUNARY0_OPMVV_rs1_vmsbf = {32'b010100_?_?????_00001_010_?????_1010111};
wildcard VMUNARY0_OPMVV_rs1_vmsof = {32'b010100_?_?????_00010_010_?????_1010111};
wildcard VMUNARY0_OPMVV_rs1_vmsif = {32'b010100_?_?????_00011_010_?????_1010111};
wildcard VMUNARY0_OPMVV_rs1_viota = {32'b010100_?_?????_10000_010_?????_1010111};
wildcard VMUNARY0_OPMVV_rs1_vid = {32'b010100_?_?????_10001_010_?????_1010111};
